* Diode Clipper Circuit
R1 n3 n2  1K
R2 n2 n1  3.3K
R3 0 n2  3.3K
R4 0 n4  5.6K

C1 n4 n2  0.47U

Vin n3 0 DC 1
Vcc1 n1 0 DC 5

D1 n2  n1 D1N3940
D2 0  n2 D1N3940
.MODEL D1N3940 D(
    + IS=4E-10 RS=.0 N=1.48 TT=8E-7
    + CJO=1.95E-11 VJ=.4 M=.38 EG=1.36
    + XTI=-8 KF=0 AF=1 FC=.9
    + BV=600 IBV=1E-4)
* RS should be 0.105. Change it when Rs is implemented in PyHBSim

.DC VIN -10 15 1
.PRINT DC file=circuit3.prn V(n3) V(n2) V(n4)

.END
